/*
*----------------------------------------------------------------------
* Module:   adder
* Function: Full Adder implemented using logic gates.
* Author:   Bibek Bhattarai
* Date:     Nov 2025
*----------------------------------------------------------------------
*/


module adder (
   input logic a,
   input logic b,
   input logic c_in,
   output logic s,
   output logic c_out
);

   assign s = a ^ b ^ c_in;
   assign c_out = (a & b) | (b & c_in) | (a & c_in);
endmodule
