module arithmetic_unit (
   logic s[3:0],
   logic a[3:0],
   logic b[3:0],
   logic f[3:0]
)

endmodule